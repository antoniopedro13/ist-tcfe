*
*NGSPICE simulation script lab1
*Group 1
*


.options savecurrents

*supply voltage

* input voltage source
Va 4 5 5.22319986769
R1 4 3 1.00676538952k
R2 2 3 2.03303206695k
R3 3 7 3.03391315228k
R4 7 5 4.00312807132k
R5 7 1 3.13101052342k
R6 5 8 2.0938993245k
R7 6 0 1.01774389701k
Id 0 1 1.03536137445m
Gb 1 2 (3,7) 7.2727641018m
Hc 7 0 Ve 8.17006533463k
Ve 8 6 0

.model group 1

.control

op

echo "**************************"
echo "Operating point"
echo "**************************"

echo "op_TAB"
print all
echo "op_END"

.endc

.end
